module ROM0 (
    input logic [3:0] addRom,
    output logic [31:0] dataRom
);
    logic [31:0] rom [15:0];

    initial begin
      rom[0]  = 32'b00000000000000000000000000000000;
		rom[1]  = 32'b00000000000000000000000000000000;
		rom[2]  = 32'b00000000000000000000000000000000;
		rom[3]  = 32'b00000000000000000000000000000000;
		rom[4]  = 32'b00000000000000000000000000000000;
		rom[5]  = 32'b00000000000001110000000000000000;
		rom[6]  = 32'b00000000000111111111111100000000;
		rom[7]  = 32'b00000000001111111111111100000000;
		rom[8]  = 32'b00000000001111111111111100000000;
		rom[9]  = 32'b00000000000111111111111100000000;
		rom[10] = 32'b00000000000001110000000000000000;
		rom[11] = 32'b00000000000000000000000000000000;
		rom[12] = 32'b00000000000000000000000000000000;
		rom[13] = 32'b00000000000000000000000000000000;
		rom[14] = 32'b00000000000000000000000000000000;
		rom[15] = 32'b00000000000000000000000000000000;
    end

    assign dataRom = rom[addRom];
	 
endmodule


module ROM1 (
    input logic [3:0] addRom,
    output logic [31:0] dataRom
);
    logic [31:0] rom [15:0];

    initial begin
        rom[0]  = 32'b00000000000000000000000000000000;
        rom[1]  = 32'b00000000000000000000000000000000;
        rom[2]  = 32'b00000000000000000000000000000000;
        rom[3]  = 32'b00000000000000000000000000000000;
        rom[4]  = 32'b00000000000000000000000000000000;
        rom[5]  = 32'b00000000000000111000000000000000;
        rom[6]  = 32'b00000011111111111110000000000000;
        rom[7]  = 32'b00000011111111111111100000000000;
        rom[8]  = 32'b00000011111111111111100000000000;
        rom[9]  = 32'b00000011111111111110000000000000;
        rom[10] = 32'b00000000000000111000000000000000;
        rom[11] = 32'b00000000000000000000000000000000;
        rom[12] = 32'b00000000000000000000000000000000;
        rom[13] = 32'b00000000000000000000000000000000;
        rom[14] = 32'b00000000000000000000000000000000;
        rom[15] = 32'b00000000000000000000000000000000;
    end

    assign dataRom = rom[addRom];
endmodule



module ROM2 (
    input logic [4:0] addRom, // Cambié a 4:0 para un rango de 0-23
    output logic [39:0] dataRom
); 
	logic [39:0] rom [23:0]; // Asegúrate de que sean 40 bits por ubicación
	initial begin
rom[0]  = 40'b0000000000000000000000110000000000000000;
rom[1]  = 40'b1111111111111111111111111111111111111111;
rom[2]  = 40'b1111111111111111111111111111111111111111;
rom[3]  = 40'b0000000000000000000000000000000000000110;
rom[4]  = 40'b0000000000000000000000000000000000001111;
rom[5]  = 40'b0000000000000111110000000000000000001111;
rom[6]  = 40'b0000000000001111111000000000000000011110;
rom[7]  = 40'b0000000000011111111100000000000000111110;
rom[8]  = 40'b0000000011111111111111111111111111111111;
rom[9]  = 40'b0000011111111111111111111111111111111111;
rom[10] = 40'b0000111000011111111111111111111111111111;
rom[11] = 40'b0001100000001111111111111111111110011110;
rom[12] = 40'b0001100001111111111111111110000000011100;
rom[13] = 40'b0011000001111111111111110000000000001100;
rom[14] = 40'b0110000001111111111110000000000000000000;
rom[15] = 40'b0100000001111111111111000000000000000000;
rom[16] = 40'b1111111111111111111111000000000000000000;
rom[17] = 40'b1111111111111111111111000000000000000000;
rom[18] = 40'b0111111111111111111110000000000000000000;
rom[19] = 40'b0111111111111111111100000000000000000000;
rom[20] = 40'b0001111111111111111000000000000000000000;
rom[21] = 40'b1000011000000000000000000000000000000000;
rom[22] = 40'b1110011000000000000000000000000000000000;
rom[23] = 40'b0111111111111111111000000000000000000000;
    end
   

    assign dataRom = rom[addRom];
endmodule


module ROM3 (
    input logic [4:0] addRom, // Cambié a 4:0 para un rango de 0-23
    output logic [39:0] dataRom
);
    logic [39:0] rom [23:0]; // Asegúrate de que sean 40 bits por ubicación

   

	 initial begin
        rom[0]  = 40'b0000000000000000000000011000000000000000;
        rom[1]  = 40'b0000000001111111111111111111111111111111;
        rom[2]  = 40'b0000000001111111111111111111111111111111;
        rom[3]  = 40'b0110000000000000000000000000000000000000;
        rom[4]  = 40'b1111000000000000000000000000000000000000;
        rom[5]  = 40'b1111000000000000000001111100000000000000;
        rom[6]  = 40'b0111100000000000000011111100000000000000;
        rom[7]  = 40'b0111110000000000000111111110000000000000;
        rom[8]  = 40'b1111111111111111111111111111110000000000;
        rom[9]  = 40'b1111111111111111111111111111111110000000;
        rom[10] = 40'b1111111111111111111111111111000011100000;
        rom[11] = 40'b0111110011111111111111111111000000110000;
        rom[12] = 40'b0011100000001111111111111111100000011000;
        rom[13] = 40'b0011000000000011111111111111100000001100;
        rom[14] = 40'b0000000000000001111111111111100000000110;
        rom[15] = 40'b0000000000000000111111111111110000000010;
        rom[16] = 40'b0000000000000000011111111111111111111111;
        rom[17] = 40'b0000000000000000011111111111111111111111;
        rom[18] = 40'b0000000000000000001111111111111111111110;
        rom[19] = 40'b0000000000000000000111111111111111111110;
        rom[20] = 40'b0000000000000000000011111111111111111000;
        rom[21] = 40'b0000000000000000000000000001000001100001;
        rom[22] = 40'b0000000000000000000000000001000001100111;
        rom[23] = 40'b0000000000000000000111111111111111111110;
    end

    assign dataRom = rom[addRom];
endmodule

